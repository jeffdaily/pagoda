netcdf fill {

dimensions:
    dim1 = 10;

variables:
    float   first(dim1);
    int     second(dim1);
    double  third(dim1);

    float   first:_FillValue = 1.0;
    char    second:missing_value = "2";

data:
    first   = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9;
    second  = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9;
    third   = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9;
}
