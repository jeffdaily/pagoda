netcdf test_pgecat1 {
dimensions:
	two = 2 ;
	three = 3 ;
	four = 4 ;
	five = 5 ;
	time = UNLIMITED ; // (0 currently)
variables:
	float two(two) ;
		two:name = "coordinate var for two" ;
	float three(three) ;
		three:name = "coordinate var for three" ;
	float four(four) ;
		four:name = "coordinate var for four" ;
	float five(five) ;
		five:name = "coordinate var for five" ;
	double a(two, three, four, five) ;
	double b(five, four, three, two) ;
	int c(three, five) ;
data:

 two = 1, 2 ;

 three = 1, 2, 3 ;

 four = 1, 2, 3, 4 ;

 five = 1, 2, 3, 4, 5 ;

 a =
  0, 1, 2, 3, 4,
  5, 6, 7, 8, 9,
  10, 11, 12, 13, 14,
  15, 16, 17, 18, 19,
  20, 21, 22, 23, 24,
  25, 26, 27, 28, 29,
  30, 31, 32, 33, 34,
  35, 36, 37, 38, 39,
  40, 41, 42, 43, 44,
  45, 46, 47, 48, 49,
  50, 51, 52, 53, 54,
  55, 56, 57, 58, 59,
  60, 61, 62, 63, 64,
  65, 66, 67, 68, 69,
  70, 71, 72, 73, 74,
  75, 76, 77, 78, 79,
  80, 81, 82, 83, 84,
  85, 86, 87, 88, 89,
  90, 91, 92, 93, 94,
  95, 96, 97, 98, 99,
  100, 101, 102, 103, 104,
  105, 106, 107, 108, 109,
  110, 111, 112, 113, 114,
  115, 116, 117, 118, 119 ;

 b =
  0, 1,
  2, 3,
  4, 5,
  6, 7,
  8, 9,
  10, 11,
  12, 13,
  14, 15,
  16, 17,
  18, 19,
  20, 21,
  22, 23,
  24, 25,
  26, 27,
  28, 29,
  30, 31,
  32, 33,
  34, 35,
  36, 37,
  38, 39,
  40, 41,
  42, 43,
  44, 45,
  46, 47,
  48, 49,
  50, 51,
  52, 53,
  54, 55,
  56, 57,
  58, 59,
  60, 61,
  62, 63,
  64, 65,
  66, 67,
  68, 69,
  70, 71,
  72, 73,
  74, 75,
  76, 77,
  78, 79,
  80, 81,
  82, 83,
  84, 85,
  86, 87,
  88, 89,
  90, 91,
  92, 93,
  94, 95,
  96, 97,
  98, 99,
  100, 101,
  102, 103,
  104, 105,
  106, 107,
  108, 109,
  110, 111,
  112, 113,
  114, 115,
  116, 117,
  118, 119 ;

 c =
  0, 1, 2, 3, 4,
  5, 6, 7, 8, 9,
  10, 11, 12, 13, 14 ;
}
